// DE10_NANO_QSYS.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module DE10_NANO_QSYS (
		output wire       adc_ltc2308_conduit_end_convst, // adc_ltc2308_conduit_end.convst
		output wire       adc_ltc2308_conduit_end_sck,    //                        .sck
		output wire       adc_ltc2308_conduit_end_sdi,    //                        .sdi
		input  wire       adc_ltc2308_conduit_end_sdo,    //                        .sdo
		input  wire       adc_ltc2308_conduit_end_dec,    //                        .dec
		input  wire       clk_clk,                        //                     clk.clk
		input  wire       i2c_dac_serial_sda_in,          //          i2c_dac_serial.sda_in
		input  wire       i2c_dac_serial_scl_in,          //                        .scl_in
		output wire       i2c_dac_serial_sda_oe,          //                        .sda_oe
		output wire       i2c_dac_serial_scl_oe,          //                        .scl_oe
		output wire       pll_sys_locked_export,          //          pll_sys_locked.export
		output wire       pll_sys_outclk2_clk,            //         pll_sys_outclk2.clk
		input  wire       reset_reset_n,                  //                   reset.reset_n
		input  wire [9:0] sw_external_connection_export   //  sw_external_connection.export
	);

	wire         pll_sys_outclk0_clk;                                                           // pll_sys:outclk_0 -> [adc_ltc2308:slave_clk, i2c_dac:clk, irq_mapper:clk, jtag_uart:clk, mm_interconnect_0:pll_sys_outclk0_clk, nios2_qsys:clk, onchip_memory2:clk, rst_controller_001:clk, rst_controller_002:clk, sw:clk, sysid_qsys:clock, timer_0:clk]
	wire         pll_sys_outclk1_clk;                                                           // pll_sys:outclk_1 -> [adc_ltc2308:adc_clk, rst_controller:clk]
	wire  [31:0] nios2_qsys_custom_instruction_master_multi_dataa;                              // nios2_qsys:A_ci_multi_dataa -> nios2_qsys_custom_instruction_master_translator:ci_slave_multi_dataa
	wire         nios2_qsys_custom_instruction_master_multi_writerc;                            // nios2_qsys:A_ci_multi_writerc -> nios2_qsys_custom_instruction_master_translator:ci_slave_multi_writerc
	wire  [31:0] nios2_qsys_custom_instruction_master_multi_result;                             // nios2_qsys_custom_instruction_master_translator:ci_slave_multi_result -> nios2_qsys:A_ci_multi_result
	wire         nios2_qsys_custom_instruction_master_clk;                                      // nios2_qsys:A_ci_multi_clock -> nios2_qsys_custom_instruction_master_translator:ci_slave_multi_clk
	wire  [31:0] nios2_qsys_custom_instruction_master_multi_datab;                              // nios2_qsys:A_ci_multi_datab -> nios2_qsys_custom_instruction_master_translator:ci_slave_multi_datab
	wire         nios2_qsys_custom_instruction_master_start;                                    // nios2_qsys:A_ci_multi_start -> nios2_qsys_custom_instruction_master_translator:ci_slave_multi_start
	wire   [4:0] nios2_qsys_custom_instruction_master_multi_b;                                  // nios2_qsys:A_ci_multi_b -> nios2_qsys_custom_instruction_master_translator:ci_slave_multi_b
	wire   [4:0] nios2_qsys_custom_instruction_master_multi_c;                                  // nios2_qsys:A_ci_multi_c -> nios2_qsys_custom_instruction_master_translator:ci_slave_multi_c
	wire         nios2_qsys_custom_instruction_master_reset_req;                                // nios2_qsys:A_ci_multi_reset_req -> nios2_qsys_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire         nios2_qsys_custom_instruction_master_done;                                     // nios2_qsys_custom_instruction_master_translator:ci_slave_multi_done -> nios2_qsys:A_ci_multi_done
	wire   [4:0] nios2_qsys_custom_instruction_master_multi_a;                                  // nios2_qsys:A_ci_multi_a -> nios2_qsys_custom_instruction_master_translator:ci_slave_multi_a
	wire         nios2_qsys_custom_instruction_master_clk_en;                                   // nios2_qsys:A_ci_multi_clk_en -> nios2_qsys_custom_instruction_master_translator:ci_slave_multi_clken
	wire         nios2_qsys_custom_instruction_master_reset;                                    // nios2_qsys:A_ci_multi_reset -> nios2_qsys_custom_instruction_master_translator:ci_slave_multi_reset
	wire         nios2_qsys_custom_instruction_master_multi_readrb;                             // nios2_qsys:A_ci_multi_readrb -> nios2_qsys_custom_instruction_master_translator:ci_slave_multi_readrb
	wire         nios2_qsys_custom_instruction_master_multi_readra;                             // nios2_qsys:A_ci_multi_readra -> nios2_qsys_custom_instruction_master_translator:ci_slave_multi_readra
	wire   [7:0] nios2_qsys_custom_instruction_master_multi_n;                                  // nios2_qsys:A_ci_multi_n -> nios2_qsys_custom_instruction_master_translator:ci_slave_multi_n
	wire         nios2_qsys_custom_instruction_master_translator_multi_ci_master_readra;        // nios2_qsys_custom_instruction_master_translator:multi_ci_master_readra -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire   [4:0] nios2_qsys_custom_instruction_master_translator_multi_ci_master_a;             // nios2_qsys_custom_instruction_master_translator:multi_ci_master_a -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_a
	wire   [4:0] nios2_qsys_custom_instruction_master_translator_multi_ci_master_b;             // nios2_qsys_custom_instruction_master_translator:multi_ci_master_b -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_b
	wire         nios2_qsys_custom_instruction_master_translator_multi_ci_master_clk;           // nios2_qsys_custom_instruction_master_translator:multi_ci_master_clk -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         nios2_qsys_custom_instruction_master_translator_multi_ci_master_readrb;        // nios2_qsys_custom_instruction_master_translator:multi_ci_master_readrb -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire   [4:0] nios2_qsys_custom_instruction_master_translator_multi_ci_master_c;             // nios2_qsys_custom_instruction_master_translator:multi_ci_master_c -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_c
	wire         nios2_qsys_custom_instruction_master_translator_multi_ci_master_start;         // nios2_qsys_custom_instruction_master_translator:multi_ci_master_start -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_start
	wire         nios2_qsys_custom_instruction_master_translator_multi_ci_master_reset_req;     // nios2_qsys_custom_instruction_master_translator:multi_ci_master_reset_req -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         nios2_qsys_custom_instruction_master_translator_multi_ci_master_done;          // nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_done -> nios2_qsys_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] nios2_qsys_custom_instruction_master_translator_multi_ci_master_n;             // nios2_qsys_custom_instruction_master_translator:multi_ci_master_n -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_n
	wire  [31:0] nios2_qsys_custom_instruction_master_translator_multi_ci_master_result;        // nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_result -> nios2_qsys_custom_instruction_master_translator:multi_ci_master_result
	wire         nios2_qsys_custom_instruction_master_translator_multi_ci_master_clk_en;        // nios2_qsys_custom_instruction_master_translator:multi_ci_master_clken -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire  [31:0] nios2_qsys_custom_instruction_master_translator_multi_ci_master_datab;         // nios2_qsys_custom_instruction_master_translator:multi_ci_master_datab -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire  [31:0] nios2_qsys_custom_instruction_master_translator_multi_ci_master_dataa;         // nios2_qsys_custom_instruction_master_translator:multi_ci_master_dataa -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         nios2_qsys_custom_instruction_master_translator_multi_ci_master_reset;         // nios2_qsys_custom_instruction_master_translator:multi_ci_master_reset -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire         nios2_qsys_custom_instruction_master_translator_multi_ci_master_writerc;       // nios2_qsys_custom_instruction_master_translator:multi_ci_master_writerc -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_readra;         // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_readra -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire   [4:0] nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_a;              // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_a -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [4:0] nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_b;              // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_b -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire         nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_readrb;         // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_readrb -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire   [4:0] nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_c;              // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_c -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_clk;            // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_clk -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire  [31:0] nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_ipending;       // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_ipending -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_start;          // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_start -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire         nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_reset_req;      // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_done;           // nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_done -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_done
	wire   [7:0] nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_n;              // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_n -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire  [31:0] nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_result;         // nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_result -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_result
	wire         nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_estatus;        // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_estatus -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire         nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_clk_en;         // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_clken -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire  [31:0] nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_datab;          // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_datab -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire  [31:0] nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_dataa;          // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_dataa -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_reset;          // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_reset -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire         nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_writerc;        // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_writerc -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_result; // recon_pipe_1_0:dac_out -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_clk;    // nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_master_clk -> recon_pipe_1_0:clk
	wire         nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_clk_en; // nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_master_clken -> recon_pipe_1_0:clk_en
	wire  [31:0] nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_dataa;  // nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> recon_pipe_1_0:adc_in
	wire         nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_start;  // nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_master_start -> recon_pipe_1_0:start
	wire         nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_reset;  // nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_master_reset -> recon_pipe_1_0:reset
	wire         nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_done;   // recon_pipe_1_0:valid_out -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire         nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_readra;         // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master1_readra -> nios2_qsys_custom_instruction_master_multi_slave_translator1:ci_slave_readra
	wire   [4:0] nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_a;              // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master1_a -> nios2_qsys_custom_instruction_master_multi_slave_translator1:ci_slave_a
	wire   [4:0] nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_b;              // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master1_b -> nios2_qsys_custom_instruction_master_multi_slave_translator1:ci_slave_b
	wire         nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_readrb;         // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master1_readrb -> nios2_qsys_custom_instruction_master_multi_slave_translator1:ci_slave_readrb
	wire   [4:0] nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_c;              // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master1_c -> nios2_qsys_custom_instruction_master_multi_slave_translator1:ci_slave_c
	wire         nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_clk;            // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master1_clk -> nios2_qsys_custom_instruction_master_multi_slave_translator1:ci_slave_clk
	wire  [31:0] nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_ipending;       // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master1_ipending -> nios2_qsys_custom_instruction_master_multi_slave_translator1:ci_slave_ipending
	wire         nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_start;          // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master1_start -> nios2_qsys_custom_instruction_master_multi_slave_translator1:ci_slave_start
	wire         nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_reset_req;      // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master1_reset_req -> nios2_qsys_custom_instruction_master_multi_slave_translator1:ci_slave_reset_req
	wire         nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_done;           // nios2_qsys_custom_instruction_master_multi_slave_translator1:ci_slave_done -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_master1_done
	wire   [7:0] nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_n;              // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master1_n -> nios2_qsys_custom_instruction_master_multi_slave_translator1:ci_slave_n
	wire  [31:0] nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_result;         // nios2_qsys_custom_instruction_master_multi_slave_translator1:ci_slave_result -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_master1_result
	wire         nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_estatus;        // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master1_estatus -> nios2_qsys_custom_instruction_master_multi_slave_translator1:ci_slave_estatus
	wire         nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_clk_en;         // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master1_clken -> nios2_qsys_custom_instruction_master_multi_slave_translator1:ci_slave_clken
	wire  [31:0] nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_datab;          // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master1_datab -> nios2_qsys_custom_instruction_master_multi_slave_translator1:ci_slave_datab
	wire  [31:0] nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_dataa;          // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master1_dataa -> nios2_qsys_custom_instruction_master_multi_slave_translator1:ci_slave_dataa
	wire         nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_reset;          // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master1_reset -> nios2_qsys_custom_instruction_master_multi_slave_translator1:ci_slave_reset
	wire         nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_writerc;        // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master1_writerc -> nios2_qsys_custom_instruction_master_multi_slave_translator1:ci_slave_writerc
	wire  [31:0] nios2_qsys_custom_instruction_master_multi_slave_translator1_ci_master_result; // recon_pipe_n_0:dac_out -> nios2_qsys_custom_instruction_master_multi_slave_translator1:ci_master_result
	wire         nios2_qsys_custom_instruction_master_multi_slave_translator1_ci_master_clk;    // nios2_qsys_custom_instruction_master_multi_slave_translator1:ci_master_clk -> recon_pipe_n_0:clk
	wire         nios2_qsys_custom_instruction_master_multi_slave_translator1_ci_master_clk_en; // nios2_qsys_custom_instruction_master_multi_slave_translator1:ci_master_clken -> recon_pipe_n_0:clk_en
	wire  [31:0] nios2_qsys_custom_instruction_master_multi_slave_translator1_ci_master_datab;  // nios2_qsys_custom_instruction_master_multi_slave_translator1:ci_master_datab -> recon_pipe_n_0:n
	wire  [31:0] nios2_qsys_custom_instruction_master_multi_slave_translator1_ci_master_dataa;  // nios2_qsys_custom_instruction_master_multi_slave_translator1:ci_master_dataa -> recon_pipe_n_0:adc_in
	wire         nios2_qsys_custom_instruction_master_multi_slave_translator1_ci_master_start;  // nios2_qsys_custom_instruction_master_multi_slave_translator1:ci_master_start -> recon_pipe_n_0:start
	wire         nios2_qsys_custom_instruction_master_multi_slave_translator1_ci_master_reset;  // nios2_qsys_custom_instruction_master_multi_slave_translator1:ci_master_reset -> recon_pipe_n_0:reset
	wire         nios2_qsys_custom_instruction_master_multi_slave_translator1_ci_master_done;   // recon_pipe_n_0:valid_out -> nios2_qsys_custom_instruction_master_multi_slave_translator1:ci_master_done
	wire  [31:0] nios2_qsys_data_master_readdata;                                               // mm_interconnect_0:nios2_qsys_data_master_readdata -> nios2_qsys:d_readdata
	wire         nios2_qsys_data_master_waitrequest;                                            // mm_interconnect_0:nios2_qsys_data_master_waitrequest -> nios2_qsys:d_waitrequest
	wire         nios2_qsys_data_master_debugaccess;                                            // nios2_qsys:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_data_master_debugaccess
	wire  [19:0] nios2_qsys_data_master_address;                                                // nios2_qsys:d_address -> mm_interconnect_0:nios2_qsys_data_master_address
	wire   [3:0] nios2_qsys_data_master_byteenable;                                             // nios2_qsys:d_byteenable -> mm_interconnect_0:nios2_qsys_data_master_byteenable
	wire         nios2_qsys_data_master_read;                                                   // nios2_qsys:d_read -> mm_interconnect_0:nios2_qsys_data_master_read
	wire         nios2_qsys_data_master_readdatavalid;                                          // mm_interconnect_0:nios2_qsys_data_master_readdatavalid -> nios2_qsys:d_readdatavalid
	wire         nios2_qsys_data_master_write;                                                  // nios2_qsys:d_write -> mm_interconnect_0:nios2_qsys_data_master_write
	wire  [31:0] nios2_qsys_data_master_writedata;                                              // nios2_qsys:d_writedata -> mm_interconnect_0:nios2_qsys_data_master_writedata
	wire  [31:0] nios2_qsys_instruction_master_readdata;                                        // mm_interconnect_0:nios2_qsys_instruction_master_readdata -> nios2_qsys:i_readdata
	wire         nios2_qsys_instruction_master_waitrequest;                                     // mm_interconnect_0:nios2_qsys_instruction_master_waitrequest -> nios2_qsys:i_waitrequest
	wire  [19:0] nios2_qsys_instruction_master_address;                                         // nios2_qsys:i_address -> mm_interconnect_0:nios2_qsys_instruction_master_address
	wire         nios2_qsys_instruction_master_read;                                            // nios2_qsys:i_read -> mm_interconnect_0:nios2_qsys_instruction_master_read
	wire         nios2_qsys_instruction_master_readdatavalid;                                   // mm_interconnect_0:nios2_qsys_instruction_master_readdatavalid -> nios2_qsys:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;                      // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;                        // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;                     // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                            // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;                       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;                           // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;                            // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire  [31:0] mm_interconnect_0_i2c_dac_csr_readdata;                                        // i2c_dac:readdata -> mm_interconnect_0:i2c_dac_csr_readdata
	wire   [3:0] mm_interconnect_0_i2c_dac_csr_address;                                         // mm_interconnect_0:i2c_dac_csr_address -> i2c_dac:addr
	wire         mm_interconnect_0_i2c_dac_csr_read;                                            // mm_interconnect_0:i2c_dac_csr_read -> i2c_dac:read
	wire         mm_interconnect_0_i2c_dac_csr_write;                                           // mm_interconnect_0:i2c_dac_csr_write -> i2c_dac:write
	wire  [31:0] mm_interconnect_0_i2c_dac_csr_writedata;                                       // mm_interconnect_0:i2c_dac_csr_writedata -> i2c_dac:writedata
	wire  [31:0] mm_interconnect_0_nios2_qsys_debug_mem_slave_readdata;                         // nios2_qsys:debug_mem_slave_readdata -> mm_interconnect_0:nios2_qsys_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_qsys_debug_mem_slave_waitrequest;                      // nios2_qsys:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_qsys_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_qsys_debug_mem_slave_debugaccess;                      // mm_interconnect_0:nios2_qsys_debug_mem_slave_debugaccess -> nios2_qsys:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_qsys_debug_mem_slave_address;                          // mm_interconnect_0:nios2_qsys_debug_mem_slave_address -> nios2_qsys:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_qsys_debug_mem_slave_read;                             // mm_interconnect_0:nios2_qsys_debug_mem_slave_read -> nios2_qsys:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_qsys_debug_mem_slave_byteenable;                       // mm_interconnect_0:nios2_qsys_debug_mem_slave_byteenable -> nios2_qsys:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_qsys_debug_mem_slave_write;                            // mm_interconnect_0:nios2_qsys_debug_mem_slave_write -> nios2_qsys:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_qsys_debug_mem_slave_writedata;                        // mm_interconnect_0:nios2_qsys_debug_mem_slave_writedata -> nios2_qsys:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_s1_chipselect;                                // mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_readdata;                                  // onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	wire  [15:0] mm_interconnect_0_onchip_memory2_s1_address;                                   // mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_s1_byteenable;                                // mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	wire         mm_interconnect_0_onchip_memory2_s1_write;                                     // mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_writedata;                                 // mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	wire         mm_interconnect_0_onchip_memory2_s1_clken;                                     // mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	wire         mm_interconnect_0_sw_s1_chipselect;                                            // mm_interconnect_0:sw_s1_chipselect -> sw:chipselect
	wire  [31:0] mm_interconnect_0_sw_s1_readdata;                                              // sw:readdata -> mm_interconnect_0:sw_s1_readdata
	wire   [1:0] mm_interconnect_0_sw_s1_address;                                               // mm_interconnect_0:sw_s1_address -> sw:address
	wire         mm_interconnect_0_sw_s1_write;                                                 // mm_interconnect_0:sw_s1_write -> sw:write_n
	wire  [31:0] mm_interconnect_0_sw_s1_writedata;                                             // mm_interconnect_0:sw_s1_writedata -> sw:writedata
	wire         mm_interconnect_0_timer_0_s1_chipselect;                                       // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                                         // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                                          // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                                            // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                                        // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_adc_ltc2308_slave_chipselect;                                // mm_interconnect_0:adc_ltc2308_slave_chipselect -> adc_ltc2308:slave_chipselect_n
	wire  [15:0] mm_interconnect_0_adc_ltc2308_slave_readdata;                                  // adc_ltc2308:slave_readdata -> mm_interconnect_0:adc_ltc2308_slave_readdata
	wire   [0:0] mm_interconnect_0_adc_ltc2308_slave_address;                                   // mm_interconnect_0:adc_ltc2308_slave_address -> adc_ltc2308:slave_addr
	wire         mm_interconnect_0_adc_ltc2308_slave_read;                                      // mm_interconnect_0:adc_ltc2308_slave_read -> adc_ltc2308:slave_read_n
	wire         mm_interconnect_0_adc_ltc2308_slave_write;                                     // mm_interconnect_0:adc_ltc2308_slave_write -> adc_ltc2308:slave_wrtie_n
	wire  [15:0] mm_interconnect_0_adc_ltc2308_slave_writedata;                                 // mm_interconnect_0:adc_ltc2308_slave_writedata -> adc_ltc2308:slave_wriredata
	wire         irq_mapper_receiver0_irq;                                                      // i2c_dac:intr -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                      // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                      // sw:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                                      // timer_0:irq -> irq_mapper:receiver3_irq
	wire  [31:0] nios2_qsys_irq_irq;                                                            // irq_mapper:sender_irq -> nios2_qsys:irq
	wire         rst_controller_reset_out_reset;                                                // rst_controller:reset_out -> adc_ltc2308:slave_reset_n
	wire         rst_controller_001_reset_out_reset;                                            // rst_controller_001:reset_out -> [i2c_dac:rst_n, jtag_uart:rst_n, mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset, onchip_memory2:reset, rst_translator:in_reset, sw:reset_n, sysid_qsys:reset_n, timer_0:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                                        // rst_controller_001:reset_req -> [onchip_memory2:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_002_reset_out_reset;                                            // rst_controller_002:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_qsys_reset_reset_bridge_in_reset_reset, nios2_qsys:reset_n]
	wire         rst_controller_002_reset_out_reset_req;                                        // rst_controller_002:reset_req -> [nios2_qsys:reset_req, rst_translator_001:reset_req_in]
	wire         nios2_qsys_debug_reset_request_reset;                                          // nios2_qsys:debug_reset_request -> rst_controller_002:reset_in1

	adc_ltc2308_fifo adc_ltc2308 (
		.slave_chipselect_n (~mm_interconnect_0_adc_ltc2308_slave_chipselect), //          slave.chipselect_n
		.slave_read_n       (~mm_interconnect_0_adc_ltc2308_slave_read),       //               .read_n
		.slave_readdata     (mm_interconnect_0_adc_ltc2308_slave_readdata),    //               .readdata
		.slave_addr         (mm_interconnect_0_adc_ltc2308_slave_address),     //               .address
		.slave_wrtie_n      (~mm_interconnect_0_adc_ltc2308_slave_write),      //               .write_n
		.slave_wriredata    (mm_interconnect_0_adc_ltc2308_slave_writedata),   //               .writedata
		.ADC_CONVST         (adc_ltc2308_conduit_end_convst),                  //    conduit_end.convst
		.ADC_SCK            (adc_ltc2308_conduit_end_sck),                     //               .sck
		.ADC_SDI            (adc_ltc2308_conduit_end_sdi),                     //               .sdi
		.ADC_SDO            (adc_ltc2308_conduit_end_sdo),                     //               .sdo
		.DEC                (adc_ltc2308_conduit_end_dec),                     //               .dec
		.adc_clk            (pll_sys_outclk1_clk),                             // clock_sink_adc.clk
		.slave_clk          (pll_sys_outclk0_clk),                             //     clock_sink.clk
		.slave_reset_n      (~rst_controller_reset_out_reset)                  //     reset_sink.reset_n
	);

	altera_avalon_i2c #(
		.USE_AV_ST       (0),
		.FIFO_DEPTH      (8),
		.FIFO_DEPTH_LOG2 (3)
	) i2c_dac (
		.clk       (pll_sys_outclk0_clk),                     //            clock.clk
		.rst_n     (~rst_controller_001_reset_out_reset),     //       reset_sink.reset_n
		.intr      (irq_mapper_receiver0_irq),                // interrupt_sender.irq
		.addr      (mm_interconnect_0_i2c_dac_csr_address),   //              csr.address
		.read      (mm_interconnect_0_i2c_dac_csr_read),      //                 .read
		.write     (mm_interconnect_0_i2c_dac_csr_write),     //                 .write
		.writedata (mm_interconnect_0_i2c_dac_csr_writedata), //                 .writedata
		.readdata  (mm_interconnect_0_i2c_dac_csr_readdata),  //                 .readdata
		.sda_in    (i2c_dac_serial_sda_in),                   //       i2c_serial.sda_in
		.scl_in    (i2c_dac_serial_scl_in),                   //                 .scl_in
		.sda_oe    (i2c_dac_serial_sda_oe),                   //                 .sda_oe
		.scl_oe    (i2c_dac_serial_scl_oe),                   //                 .scl_oe
		.src_data  (),                                        //      (terminated)
		.src_valid (),                                        //      (terminated)
		.src_ready (1'b0),                                    //      (terminated)
		.snk_data  (16'b0000000000000000),                    //      (terminated)
		.snk_valid (1'b0),                                    //      (terminated)
		.snk_ready ()                                         //      (terminated)
	);

	DE10_NANO_QSYS_jtag_uart jtag_uart (
		.clk            (pll_sys_outclk0_clk),                                       //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	DE10_NANO_QSYS_nios2_qsys nios2_qsys (
		.clk                                 (pll_sys_outclk0_clk),                                      //                       clk.clk
		.reset_n                             (~rst_controller_002_reset_out_reset),                      //                     reset.reset_n
		.reset_req                           (rst_controller_002_reset_out_reset_req),                   //                          .reset_req
		.d_address                           (nios2_qsys_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_qsys_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_qsys_data_master_read),                              //                          .read
		.d_readdata                          (nios2_qsys_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_qsys_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_qsys_data_master_write),                             //                          .write
		.d_writedata                         (nios2_qsys_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_qsys_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_qsys_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_qsys_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_qsys_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_qsys_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_qsys_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_qsys_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_qsys_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_qsys_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_qsys_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_qsys_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_qsys_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_qsys_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_qsys_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_qsys_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_qsys_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_qsys_debug_mem_slave_writedata),   //                          .writedata
		.A_ci_multi_done                     (nios2_qsys_custom_instruction_master_done),                // custom_instruction_master.done
		.A_ci_multi_result                   (nios2_qsys_custom_instruction_master_multi_result),        //                          .multi_result
		.A_ci_multi_a                        (nios2_qsys_custom_instruction_master_multi_a),             //                          .multi_a
		.A_ci_multi_b                        (nios2_qsys_custom_instruction_master_multi_b),             //                          .multi_b
		.A_ci_multi_c                        (nios2_qsys_custom_instruction_master_multi_c),             //                          .multi_c
		.A_ci_multi_clk_en                   (nios2_qsys_custom_instruction_master_clk_en),              //                          .clk_en
		.A_ci_multi_clock                    (nios2_qsys_custom_instruction_master_clk),                 //                          .clk
		.A_ci_multi_reset                    (nios2_qsys_custom_instruction_master_reset),               //                          .reset
		.A_ci_multi_reset_req                (nios2_qsys_custom_instruction_master_reset_req),           //                          .reset_req
		.A_ci_multi_dataa                    (nios2_qsys_custom_instruction_master_multi_dataa),         //                          .multi_dataa
		.A_ci_multi_datab                    (nios2_qsys_custom_instruction_master_multi_datab),         //                          .multi_datab
		.A_ci_multi_n                        (nios2_qsys_custom_instruction_master_multi_n),             //                          .multi_n
		.A_ci_multi_readra                   (nios2_qsys_custom_instruction_master_multi_readra),        //                          .multi_readra
		.A_ci_multi_readrb                   (nios2_qsys_custom_instruction_master_multi_readrb),        //                          .multi_readrb
		.A_ci_multi_start                    (nios2_qsys_custom_instruction_master_start),               //                          .start
		.A_ci_multi_writerc                  (nios2_qsys_custom_instruction_master_multi_writerc)        //                          .multi_writerc
	);

	DE10_NANO_QSYS_onchip_memory2 onchip_memory2 (
		.clk        (pll_sys_outclk0_clk),                            //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),         //       .reset_req
		.freeze     (1'b0)                                            // (terminated)
	);

	DE10_NANO_QSYS_pll_sys pll_sys (
		.refclk   (clk_clk),               //  refclk.clk
		.rst      (~reset_reset_n),        //   reset.reset
		.outclk_0 (pll_sys_outclk0_clk),   // outclk0.clk
		.outclk_1 (pll_sys_outclk1_clk),   // outclk1.clk
		.outclk_2 (pll_sys_outclk2_clk),   // outclk2.clk
		.locked   (pll_sys_locked_export)  //  locked.export
	);

	reconstruction_top_pipelined #(
		.WIDTH           (24),
		.LAMBDA          (26'b00000000010001100110011010),
		.FRACTIONAL_BITS (16),
		.WINDOW_SIZE     (100),
		.one_over_a      (6554)
	) recon_pipe_1_0 (
		.clk_en    (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), // nios_custom_instruction_slave.clk_en
		.start     (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_start),  //                              .start
		.adc_in    (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  //                              .dataa
		.valid_out (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_done),   //                              .done
		.dac_out   (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_result), //                              .result
		.clk       (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //                              .clk
		.reset     (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_reset)   //                              .reset
	);

	reconstruction_top_pipelined_n #(
		.WIDTH           (24),
		.LAMBDA          (26'b00000000010001100110011010),
		.FRACTIONAL_BITS (16),
		.WINDOW_SIZE     (100),
		.one_over_a      (6554)
	) recon_pipe_n_0 (
		.clk_en    (nios2_qsys_custom_instruction_master_multi_slave_translator1_ci_master_clk_en), // nios_custom_instruction_slave.clk_en
		.start     (nios2_qsys_custom_instruction_master_multi_slave_translator1_ci_master_start),  //                              .start
		.adc_in    (nios2_qsys_custom_instruction_master_multi_slave_translator1_ci_master_dataa),  //                              .dataa
		.n         (nios2_qsys_custom_instruction_master_multi_slave_translator1_ci_master_datab),  //                              .datab
		.valid_out (nios2_qsys_custom_instruction_master_multi_slave_translator1_ci_master_done),   //                              .done
		.dac_out   (nios2_qsys_custom_instruction_master_multi_slave_translator1_ci_master_result), //                              .result
		.clk       (nios2_qsys_custom_instruction_master_multi_slave_translator1_ci_master_clk),    //                              .clk
		.reset     (nios2_qsys_custom_instruction_master_multi_slave_translator1_ci_master_reset)   //                              .reset
	);

	DE10_NANO_QSYS_sw sw (
		.clk        (pll_sys_outclk0_clk),                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_0_sw_s1_address),     //                  s1.address
		.write_n    (~mm_interconnect_0_sw_s1_write),      //                    .write_n
		.writedata  (mm_interconnect_0_sw_s1_writedata),   //                    .writedata
		.chipselect (mm_interconnect_0_sw_s1_chipselect),  //                    .chipselect
		.readdata   (mm_interconnect_0_sw_s1_readdata),    //                    .readdata
		.in_port    (sw_external_connection_export),       // external_connection.export
		.irq        (irq_mapper_receiver2_irq)             //                 irq.irq
	);

	DE10_NANO_QSYS_sysid_qsys sysid_qsys (
		.clock    (pll_sys_outclk0_clk),                                 //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	DE10_NANO_QSYS_timer_0 timer_0 (
		.clk        (pll_sys_outclk0_clk),                     //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                 //   irq.irq
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (0)
	) nios2_qsys_custom_instruction_master_translator (
		.ci_slave_result           (),                                                                          //        ci_slave.result
		.ci_slave_multi_clk        (nios2_qsys_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (nios2_qsys_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (nios2_qsys_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (nios2_qsys_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (nios2_qsys_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (nios2_qsys_custom_instruction_master_done),                                 //                .done
		.ci_slave_multi_dataa      (nios2_qsys_custom_instruction_master_multi_dataa),                          //                .multi_dataa
		.ci_slave_multi_datab      (nios2_qsys_custom_instruction_master_multi_datab),                          //                .multi_datab
		.ci_slave_multi_result     (nios2_qsys_custom_instruction_master_multi_result),                         //                .multi_result
		.ci_slave_multi_n          (nios2_qsys_custom_instruction_master_multi_n),                              //                .multi_n
		.ci_slave_multi_readra     (nios2_qsys_custom_instruction_master_multi_readra),                         //                .multi_readra
		.ci_slave_multi_readrb     (nios2_qsys_custom_instruction_master_multi_readrb),                         //                .multi_readrb
		.ci_slave_multi_writerc    (nios2_qsys_custom_instruction_master_multi_writerc),                        //                .multi_writerc
		.ci_slave_multi_a          (nios2_qsys_custom_instruction_master_multi_a),                              //                .multi_a
		.ci_slave_multi_b          (nios2_qsys_custom_instruction_master_multi_b),                              //                .multi_b
		.ci_slave_multi_c          (nios2_qsys_custom_instruction_master_multi_c),                              //                .multi_c
		.comb_ci_master_result     (),                                                                          //  comb_ci_master.result
		.multi_ci_master_clk       (nios2_qsys_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (nios2_qsys_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (nios2_qsys_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (nios2_qsys_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (nios2_qsys_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (nios2_qsys_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (nios2_qsys_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (nios2_qsys_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (nios2_qsys_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (nios2_qsys_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (nios2_qsys_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (nios2_qsys_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (nios2_qsys_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (nios2_qsys_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (nios2_qsys_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (nios2_qsys_custom_instruction_master_translator_multi_ci_master_c),         //                .c
		.ci_slave_dataa            (32'b00000000000000000000000000000000),                                      //     (terminated)
		.ci_slave_datab            (32'b00000000000000000000000000000000),                                      //     (terminated)
		.ci_slave_n                (8'b00000000),                                                               //     (terminated)
		.ci_slave_readra           (1'b0),                                                                      //     (terminated)
		.ci_slave_readrb           (1'b0),                                                                      //     (terminated)
		.ci_slave_writerc          (1'b0),                                                                      //     (terminated)
		.ci_slave_a                (5'b00000),                                                                  //     (terminated)
		.ci_slave_b                (5'b00000),                                                                  //     (terminated)
		.ci_slave_c                (5'b00000),                                                                  //     (terminated)
		.ci_slave_ipending         (32'b00000000000000000000000000000000),                                      //     (terminated)
		.ci_slave_estatus          (1'b0),                                                                      //     (terminated)
		.comb_ci_master_dataa      (),                                                                          //     (terminated)
		.comb_ci_master_datab      (),                                                                          //     (terminated)
		.comb_ci_master_n          (),                                                                          //     (terminated)
		.comb_ci_master_readra     (),                                                                          //     (terminated)
		.comb_ci_master_readrb     (),                                                                          //     (terminated)
		.comb_ci_master_writerc    (),                                                                          //     (terminated)
		.comb_ci_master_a          (),                                                                          //     (terminated)
		.comb_ci_master_b          (),                                                                          //     (terminated)
		.comb_ci_master_c          (),                                                                          //     (terminated)
		.comb_ci_master_ipending   (),                                                                          //     (terminated)
		.comb_ci_master_estatus    ()                                                                           //     (terminated)
	);

	DE10_NANO_QSYS_nios2_qsys_custom_instruction_master_multi_xconnect nios2_qsys_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (nios2_qsys_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (nios2_qsys_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (nios2_qsys_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (nios2_qsys_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (nios2_qsys_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (nios2_qsys_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (nios2_qsys_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (nios2_qsys_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (nios2_qsys_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (nios2_qsys_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                          //           .ipending
		.ci_slave_estatus     (),                                                                          //           .estatus
		.ci_slave_clk         (nios2_qsys_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (nios2_qsys_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (nios2_qsys_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (nios2_qsys_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (nios2_qsys_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (nios2_qsys_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_done),       //           .done
		.ci_master1_dataa     (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_dataa),      // ci_master1.dataa
		.ci_master1_datab     (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_datab),      //           .datab
		.ci_master1_result    (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_result),     //           .result
		.ci_master1_n         (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_n),          //           .n
		.ci_master1_readra    (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_readra),     //           .readra
		.ci_master1_readrb    (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_readrb),     //           .readrb
		.ci_master1_writerc   (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_writerc),    //           .writerc
		.ci_master1_a         (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_a),          //           .a
		.ci_master1_b         (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_b),          //           .b
		.ci_master1_c         (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_c),          //           .c
		.ci_master1_ipending  (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_ipending),   //           .ipending
		.ci_master1_estatus   (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_estatus),    //           .estatus
		.ci_master1_clk       (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_clk),        //           .clk
		.ci_master1_reset     (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_reset),      //           .reset
		.ci_master1_clken     (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_clk_en),     //           .clk_en
		.ci_master1_reset_req (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_reset_req),  //           .reset_req
		.ci_master1_start     (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_start),      //           .start
		.ci_master1_done      (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) nios2_qsys_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_estatus),        //          .estatus
		.ci_slave_clk        (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_clk),            //          .clk
		.ci_slave_clken      (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_clk_en),         //          .clk_en
		.ci_slave_reset_req  (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_reset_req),      //          .reset_req
		.ci_slave_reset      (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_reset),          //          .reset
		.ci_slave_start      (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_start),          //          .start
		.ci_slave_done       (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_done),           //          .done
		.ci_master_dataa     (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_result    (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_result), //          .result
		.ci_master_clk       (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //          .clk
		.ci_master_clken     (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //          .reset
		.ci_master_start     (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_start),  //          .start
		.ci_master_done      (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_done),   //          .done
		.ci_master_datab     (),                                                                              // (terminated)
		.ci_master_n         (),                                                                              // (terminated)
		.ci_master_readra    (),                                                                              // (terminated)
		.ci_master_readrb    (),                                                                              // (terminated)
		.ci_master_writerc   (),                                                                              // (terminated)
		.ci_master_a         (),                                                                              // (terminated)
		.ci_master_b         (),                                                                              // (terminated)
		.ci_master_c         (),                                                                              // (terminated)
		.ci_master_ipending  (),                                                                              // (terminated)
		.ci_master_estatus   (),                                                                              // (terminated)
		.ci_master_reset_req ()                                                                               // (terminated)
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) nios2_qsys_custom_instruction_master_multi_slave_translator1 (
		.ci_slave_dataa      (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_datab),          //          .datab
		.ci_slave_result     (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_result),         //          .result
		.ci_slave_n          (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_n),              //          .n
		.ci_slave_readra     (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_readra),         //          .readra
		.ci_slave_readrb     (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_writerc),        //          .writerc
		.ci_slave_a          (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_a),              //          .a
		.ci_slave_b          (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_b),              //          .b
		.ci_slave_c          (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_c),              //          .c
		.ci_slave_ipending   (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_estatus),        //          .estatus
		.ci_slave_clk        (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_clk),            //          .clk
		.ci_slave_clken      (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_clk_en),         //          .clk_en
		.ci_slave_reset_req  (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_reset_req),      //          .reset_req
		.ci_slave_reset      (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_reset),          //          .reset
		.ci_slave_start      (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_start),          //          .start
		.ci_slave_done       (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master1_done),           //          .done
		.ci_master_dataa     (nios2_qsys_custom_instruction_master_multi_slave_translator1_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios2_qsys_custom_instruction_master_multi_slave_translator1_ci_master_datab),  //          .datab
		.ci_master_result    (nios2_qsys_custom_instruction_master_multi_slave_translator1_ci_master_result), //          .result
		.ci_master_clk       (nios2_qsys_custom_instruction_master_multi_slave_translator1_ci_master_clk),    //          .clk
		.ci_master_clken     (nios2_qsys_custom_instruction_master_multi_slave_translator1_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (nios2_qsys_custom_instruction_master_multi_slave_translator1_ci_master_reset),  //          .reset
		.ci_master_start     (nios2_qsys_custom_instruction_master_multi_slave_translator1_ci_master_start),  //          .start
		.ci_master_done      (nios2_qsys_custom_instruction_master_multi_slave_translator1_ci_master_done),   //          .done
		.ci_master_n         (),                                                                              // (terminated)
		.ci_master_readra    (),                                                                              // (terminated)
		.ci_master_readrb    (),                                                                              // (terminated)
		.ci_master_writerc   (),                                                                              // (terminated)
		.ci_master_a         (),                                                                              // (terminated)
		.ci_master_b         (),                                                                              // (terminated)
		.ci_master_c         (),                                                                              // (terminated)
		.ci_master_ipending  (),                                                                              // (terminated)
		.ci_master_estatus   (),                                                                              // (terminated)
		.ci_master_reset_req ()                                                                               // (terminated)
	);

	DE10_NANO_QSYS_mm_interconnect_0 mm_interconnect_0 (
		.pll_sys_outclk0_clk                          (pll_sys_outclk0_clk),                                       //                        pll_sys_outclk0.clk
		.jtag_uart_reset_reset_bridge_in_reset_reset  (rst_controller_001_reset_out_reset),                        //  jtag_uart_reset_reset_bridge_in_reset.reset
		.nios2_qsys_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                        // nios2_qsys_reset_reset_bridge_in_reset.reset
		.nios2_qsys_data_master_address               (nios2_qsys_data_master_address),                            //                 nios2_qsys_data_master.address
		.nios2_qsys_data_master_waitrequest           (nios2_qsys_data_master_waitrequest),                        //                                       .waitrequest
		.nios2_qsys_data_master_byteenable            (nios2_qsys_data_master_byteenable),                         //                                       .byteenable
		.nios2_qsys_data_master_read                  (nios2_qsys_data_master_read),                               //                                       .read
		.nios2_qsys_data_master_readdata              (nios2_qsys_data_master_readdata),                           //                                       .readdata
		.nios2_qsys_data_master_readdatavalid         (nios2_qsys_data_master_readdatavalid),                      //                                       .readdatavalid
		.nios2_qsys_data_master_write                 (nios2_qsys_data_master_write),                              //                                       .write
		.nios2_qsys_data_master_writedata             (nios2_qsys_data_master_writedata),                          //                                       .writedata
		.nios2_qsys_data_master_debugaccess           (nios2_qsys_data_master_debugaccess),                        //                                       .debugaccess
		.nios2_qsys_instruction_master_address        (nios2_qsys_instruction_master_address),                     //          nios2_qsys_instruction_master.address
		.nios2_qsys_instruction_master_waitrequest    (nios2_qsys_instruction_master_waitrequest),                 //                                       .waitrequest
		.nios2_qsys_instruction_master_read           (nios2_qsys_instruction_master_read),                        //                                       .read
		.nios2_qsys_instruction_master_readdata       (nios2_qsys_instruction_master_readdata),                    //                                       .readdata
		.nios2_qsys_instruction_master_readdatavalid  (nios2_qsys_instruction_master_readdatavalid),               //                                       .readdatavalid
		.adc_ltc2308_slave_address                    (mm_interconnect_0_adc_ltc2308_slave_address),               //                      adc_ltc2308_slave.address
		.adc_ltc2308_slave_write                      (mm_interconnect_0_adc_ltc2308_slave_write),                 //                                       .write
		.adc_ltc2308_slave_read                       (mm_interconnect_0_adc_ltc2308_slave_read),                  //                                       .read
		.adc_ltc2308_slave_readdata                   (mm_interconnect_0_adc_ltc2308_slave_readdata),              //                                       .readdata
		.adc_ltc2308_slave_writedata                  (mm_interconnect_0_adc_ltc2308_slave_writedata),             //                                       .writedata
		.adc_ltc2308_slave_chipselect                 (mm_interconnect_0_adc_ltc2308_slave_chipselect),            //                                       .chipselect
		.i2c_dac_csr_address                          (mm_interconnect_0_i2c_dac_csr_address),                     //                            i2c_dac_csr.address
		.i2c_dac_csr_write                            (mm_interconnect_0_i2c_dac_csr_write),                       //                                       .write
		.i2c_dac_csr_read                             (mm_interconnect_0_i2c_dac_csr_read),                        //                                       .read
		.i2c_dac_csr_readdata                         (mm_interconnect_0_i2c_dac_csr_readdata),                    //                                       .readdata
		.i2c_dac_csr_writedata                        (mm_interconnect_0_i2c_dac_csr_writedata),                   //                                       .writedata
		.jtag_uart_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //            jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                       .write
		.jtag_uart_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                       .read
		.jtag_uart_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                       .readdata
		.jtag_uart_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                       .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                       .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                       .chipselect
		.nios2_qsys_debug_mem_slave_address           (mm_interconnect_0_nios2_qsys_debug_mem_slave_address),      //             nios2_qsys_debug_mem_slave.address
		.nios2_qsys_debug_mem_slave_write             (mm_interconnect_0_nios2_qsys_debug_mem_slave_write),        //                                       .write
		.nios2_qsys_debug_mem_slave_read              (mm_interconnect_0_nios2_qsys_debug_mem_slave_read),         //                                       .read
		.nios2_qsys_debug_mem_slave_readdata          (mm_interconnect_0_nios2_qsys_debug_mem_slave_readdata),     //                                       .readdata
		.nios2_qsys_debug_mem_slave_writedata         (mm_interconnect_0_nios2_qsys_debug_mem_slave_writedata),    //                                       .writedata
		.nios2_qsys_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_qsys_debug_mem_slave_byteenable),   //                                       .byteenable
		.nios2_qsys_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_qsys_debug_mem_slave_waitrequest),  //                                       .waitrequest
		.nios2_qsys_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_qsys_debug_mem_slave_debugaccess),  //                                       .debugaccess
		.onchip_memory2_s1_address                    (mm_interconnect_0_onchip_memory2_s1_address),               //                      onchip_memory2_s1.address
		.onchip_memory2_s1_write                      (mm_interconnect_0_onchip_memory2_s1_write),                 //                                       .write
		.onchip_memory2_s1_readdata                   (mm_interconnect_0_onchip_memory2_s1_readdata),              //                                       .readdata
		.onchip_memory2_s1_writedata                  (mm_interconnect_0_onchip_memory2_s1_writedata),             //                                       .writedata
		.onchip_memory2_s1_byteenable                 (mm_interconnect_0_onchip_memory2_s1_byteenable),            //                                       .byteenable
		.onchip_memory2_s1_chipselect                 (mm_interconnect_0_onchip_memory2_s1_chipselect),            //                                       .chipselect
		.onchip_memory2_s1_clken                      (mm_interconnect_0_onchip_memory2_s1_clken),                 //                                       .clken
		.sw_s1_address                                (mm_interconnect_0_sw_s1_address),                           //                                  sw_s1.address
		.sw_s1_write                                  (mm_interconnect_0_sw_s1_write),                             //                                       .write
		.sw_s1_readdata                               (mm_interconnect_0_sw_s1_readdata),                          //                                       .readdata
		.sw_s1_writedata                              (mm_interconnect_0_sw_s1_writedata),                         //                                       .writedata
		.sw_s1_chipselect                             (mm_interconnect_0_sw_s1_chipselect),                        //                                       .chipselect
		.sysid_qsys_control_slave_address             (mm_interconnect_0_sysid_qsys_control_slave_address),        //               sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata            (mm_interconnect_0_sysid_qsys_control_slave_readdata),       //                                       .readdata
		.timer_0_s1_address                           (mm_interconnect_0_timer_0_s1_address),                      //                             timer_0_s1.address
		.timer_0_s1_write                             (mm_interconnect_0_timer_0_s1_write),                        //                                       .write
		.timer_0_s1_readdata                          (mm_interconnect_0_timer_0_s1_readdata),                     //                                       .readdata
		.timer_0_s1_writedata                         (mm_interconnect_0_timer_0_s1_writedata),                    //                                       .writedata
		.timer_0_s1_chipselect                        (mm_interconnect_0_timer_0_s1_chipselect)                    //                                       .chipselect
	);

	DE10_NANO_QSYS_irq_mapper irq_mapper (
		.clk           (pll_sys_outclk0_clk),                //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.sender_irq    (nios2_qsys_irq_irq)                  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (pll_sys_outclk1_clk),            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (pll_sys_outclk0_clk),                    //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_qsys_debug_reset_request_reset),   // reset_in1.reset
		.clk            (pll_sys_outclk0_clk),                    //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
